module Incrementer(input [12:0] a, output [12:0] out);
	assign out = a + 1;
endmodule
